// Bayley King, Bryan Kanu, Zach Hadden
// Embedded Systems final project
// Logic operations on 64-bit inputs

`timescale 1ns / 100ps

module int_log(clk, operation, opa, opb, out);
input       clk;
input       [2:0] operation; 
input       [63:0]  opa, opb;
output      [63:0]  out;      

reg         [63:0]  out_temp; 

always @ (clk) begin
    
    case (operation)
    3'b000: out_temp <= opa & opb;       // A & B
    3'b001: out_temp <= ~(opa & opb);    // ~(A & opb)
    3'b010: out_temp <= opa | opb;       // A x B
    3'b011: out_temp <= ~(opa | opb);    // ~(A | B)
    3'b100: out_temp <= opa ^ opb;       // A ^ B 
    3'b101: out_temp <= ~(opa ^ opb);    // ~(A^B)
    3'b110: out_temp <= !(opa);          // A^B
    endcase

end

assign out = out_temp;

endmodule